library verilog;
use verilog.vl_types.all;
entity eviction_write_buffer_sv_unit is
end eviction_write_buffer_sv_unit;
