library verilog;
use verilog.vl_types.all;
entity l2_detect_hit_sv_unit is
end l2_detect_hit_sv_unit;
