library verilog;
use verilog.vl_types.all;
entity if_id_state_reg_sv_unit is
end if_id_state_reg_sv_unit;
