library verilog;
use verilog.vl_types.all;
entity arb_control_sv_unit is
end arb_control_sv_unit;
