library verilog;
use verilog.vl_types.all;
entity perf_counters_sv_unit is
end perf_counters_sv_unit;
