library verilog;
use verilog.vl_types.all;
entity ex_mem_state_reg_sv_unit is
end ex_mem_state_reg_sv_unit;
