library verilog;
use verilog.vl_types.all;
entity id_ex_state_reg_sv_unit is
end id_ex_state_reg_sv_unit;
