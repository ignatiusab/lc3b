library verilog;
use verilog.vl_types.all;
entity pattern_history_table_sv_unit is
end pattern_history_table_sv_unit;
