library verilog;
use verilog.vl_types.all;
entity demux16_sv_unit is
end demux16_sv_unit;
