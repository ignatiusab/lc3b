library verilog;
use verilog.vl_types.all;
entity pmem_registers_sv_unit is
end pmem_registers_sv_unit;
