library verilog;
use verilog.vl_types.all;
entity demux2_sv_unit is
end demux2_sv_unit;
