library verilog;
use verilog.vl_types.all;
entity high_low_byte_selector_sv_unit is
end high_low_byte_selector_sv_unit;
