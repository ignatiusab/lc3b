library verilog;
use verilog.vl_types.all;
entity branch_target_buffer_sv_unit is
end branch_target_buffer_sv_unit;
