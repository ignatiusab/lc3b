library verilog;
use verilog.vl_types.all;
entity branch_predictor_sv_unit is
end branch_predictor_sv_unit;
