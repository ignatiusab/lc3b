library verilog;
use verilog.vl_types.all;
entity arb_datapath_sv_unit is
end arb_datapath_sv_unit;
