library verilog;
use verilog.vl_types.all;
entity l1_cache_sv_unit is
end l1_cache_sv_unit;
