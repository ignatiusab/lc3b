library verilog;
use verilog.vl_types.all;
entity mux8_sv_unit is
end mux8_sv_unit;
