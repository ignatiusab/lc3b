library verilog;
use verilog.vl_types.all;
entity local_branch_history_predictor_sv_unit is
end local_branch_history_predictor_sv_unit;
