library verilog;
use verilog.vl_types.all;
entity zext_high_low_byte_sv_unit is
end zext_high_low_byte_sv_unit;
