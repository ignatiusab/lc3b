library verilog;
use verilog.vl_types.all;
entity mux2_sv_unit is
end mux2_sv_unit;
