library verilog;
use verilog.vl_types.all;
entity detect_hit_sv_unit is
end detect_hit_sv_unit;
