library verilog;
use verilog.vl_types.all;
entity l2_line_builder_sv_unit is
end l2_line_builder_sv_unit;
