library verilog;
use verilog.vl_types.all;
entity line_builder_sv_unit is
end line_builder_sv_unit;
