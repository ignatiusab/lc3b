library verilog;
use verilog.vl_types.all;
entity waymux4_sv_unit is
end waymux4_sv_unit;
