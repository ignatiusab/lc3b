library verilog;
use verilog.vl_types.all;
entity global_branch_history_predictor_sv_unit is
end global_branch_history_predictor_sv_unit;
