library verilog;
use verilog.vl_types.all;
entity mmio_sv_unit is
end mmio_sv_unit;
