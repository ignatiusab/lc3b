library verilog;
use verilog.vl_types.all;
entity btb_entry_sv_unit is
end btb_entry_sv_unit;
